`timescale 1ns / 1ps

module ALUController (
    //Inputs
    input logic [1:0] ALUOp,  // 2-bit opcode field from the Controller--00: LW/SW/AUIPC; 01:Branch; 10: Rtype/Itype; 11:JAL/LUI
    input logic [6:0] Funct7,  // bits 25 to 31 of the instruction
    input logic [2:0] Funct3,  // bits 12 to 14 of the instruction
    //Output
    output logic [3:0] Operation  // operation selection for ALU
);
    always_comb
        begin
            case(ALUOp)
                2'b00:
                    if(Funct3 == 3'b010)    //LW SW
                        Operation = 4'b0100;
                    else
                        Operation = 4'b0000;
                2'b01:
                        Operation = 4'b1000;
                2'b10:
                    if(Funct3 == 3'b101)    //ADDI
                        Operation = 4'b0100;
                    else if(Funct3 == 3'b000 && Funct7 == 7'b0000000)   //ADD
                        Operation = 4'b0100;
                    else if(Funct3 == 3'b000 && Funct7 == 7'b0100000)   //SUB
                        Operation = 4'b0101;
                    else if(Funct3 == 3'b111 && Funct7 == 7'b0000000)   //AND
                        Operation = 4'b0000;
                    else if(Funct3 == 3'b110 && Funct7 == 7'b0000000)   //OR
                        Operation = 4'b0001;
                    else if(Funct3 == 3'b100 && Funct7 == 7'b0000000)   //XOR
                        Operation = 4'b0010;
                    else
                        Operation = 4'b0000;
                2'b11:
                        Operation = 4'b0000;
                default:
                        Operation = 4'b0000;
            endcase
        end

    // assign Operation[0] = ((ALUOp == 2'b10) && (Funct3 == 3'b110)) ||  // R\I-or
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0000000)) ||  // R\I->>
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0100000));  // R\I->>>

    // assign Operation[1] = (ALUOp == 2'b00) ||  // LW\SW
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0000000)) ||  // R\I-add
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0010011)) ||  // addi
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0100000));  // R\I->>>

    // assign Operation[2] =  ((ALUOp==2'b10) && (Funct3==3'b101) && (Funct7==7'b0000000)) || // R\I->>
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b101) && (Funct7 == 7'b0100000)) ||  // R\I->>>
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b000) && (Funct7 == 7'b0100000)) ||  // sub
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b001)) ||  // R\I-<<
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b010));  // R\I-<

    // assign Operation[3] = (ALUOp == 2'b01) ||  // BEQ
    //     ((ALUOp == 2'b10) && (Funct3 == 3'b010));  // R\I-<
endmodule
